library verilog;
use verilog.vl_types.all;
entity tst_dec_4x16 is
end tst_dec_4x16;
